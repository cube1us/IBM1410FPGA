-- START USER TEST BENCH DECLARATIONS

-- The user test bench declaraionts, if any, must be
-- placed AFTER the line starts with the first line of text 
-- that -- START USER TEST BENCH DECLARATIONS and ends
-- with --END .
-- This text is preserved when the IBM1410SMS applciation
-- regenerates a test bench

   -- Your test bench declarations go here

-- END USER TEST BENCH DECLARATIONS
   