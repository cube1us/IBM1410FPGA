----------------------------------------------------------------------------------
-- Company: The Computer Collection 
-- Engineer: Jay R. Jaeger   
-- 
-- Create Date: 05/02/2022 03:43:13 PM
-- Design Name: IBM1410
-- Module Name: IBM1410_MEMORY_LOADER_RECEIVER - Behavioral
-- Project Name: IBM1410 
-- Target Devices: 
-- Tool Versions: 
-- Description: This module receives data from the PC console host via module
--   IBM1410_UART_INPUT_SUBSYSTEM.  It uses that data to load memory.
--   Obviously, a real IBM 1410 did NOT have such a feature.  ;)
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IBM1410_MEMORY_LOADER_RECEIVER is
    Port ( FPGA_CLK : in STD_LOGIC;
           RESET : in STD_LOGIC;
           LOADER_FIFO_WRITE_ENABLE : in STD_LOGIC;
           LOADER_FIFO_WRITE_DATA : in STD_LOGIC_VECTOR (7 downto 0);
           IBM1410_DIRECT_MEMORY_ADDRESS: out STD_LOGIC_VECTOR(13 downto 0);
           IBM1410_LOADER_DIRECT_MEMORY_ENABLE:  out STD_LOGIC_VECTOR(3 downto 0);
           IBM1410_LOADER_DIRECT_MEMORY_WRITE_ENABLE:  out STD_LOGIC_VECTOR(3 downto 0);
           IBM1410_DIRECT_MEMORY_WRITE_DATA: out STD_LOGIC_VECTOR(7 downto 0)
    );
end IBM1410_CONSOLE_SWITCHES_RECEIVER;

architecture Behavioral of IBM1410_MEMORY_LOADER_RECEIVER is

   component ring_buffer is
      generic (
         RAM_WIDTH : natural;
         RAM_DEPTH : natural
      );
      port (
         clk : in std_logic;
         rst : in std_logic;

         -- Write port
         wr_en : in std_logic;
         wr_data : in std_logic_vector(RAM_WIDTH - 1 downto 0);

         -- Read port
         rd_en : in std_logic;
         rd_valid : out std_logic;
         rd_data : out std_logic_vector(RAM_WIDTH - 1 downto 0);

         -- Flags
         empty : out std_logic;
         empty_next : out std_logic;
         full : out std_logic;
         full_next : out std_logic;

         -- The number of elements in the FIFO
         fill_count : out integer range RAM_DEPTH - 1 downto 0
      );
   end component;
   
constant MEMORY_LOADER_FIFO_SIZE: INTEGER := 16;
constant MEMORY_LOADER_FIFO_WIDTH: INTEGER := 8;
constant MEMORY_LOADER_ADDRESS_MARK: STD_LOGIC_VECTOR(6 downto 0) := "1000000";
constant MEMORY_LOADER_END_MARK: STD_LOGIC_VECTOR(6 downto 0) := "1110000";
constant MEMORY_LOADER_DATA_0_MARK: STD_LOGIC_VECTOR(6 downto 0) := "0100000";
constant MEMORY_LOADER_DATA_1_MARK: STD_LOGIC_VECTOR(6 downto 0) := "0010000";


type loaderState_type is (
   loader_Reset, loader_WaitForChar, loader_Getchar, loader_Action,
	loader_Write, loader_WrDone);

type loaderAction_type is (loader_None, loader_Addr, loader_Data_0, loader_Data_1);
   

signal loaderState: loaderState_type := loader_Reset;
signal loaderAction: loaderAction_type := loader_None;

signal FIFO_READ_ENABLE:     STD_LOGIC := '0';
signal FIFO_READ_DATA_VALID: STD_LOGIC;
signal FIFO_READ_DATA:       STD_LOGIC_VECTOR(7 downto 0);
signal FIFO_EMPTY:           STD_LOGIC;
signal FIFO_EMPTY_NEXT:      STD_LOGIC;
signal FIFO_FULL: STD_LOGIC;        -- Not used - assumption for now is that 1410 will keep up.
signal FIFO_FULL_NEXT: STD_LOGIC;   -- Not used - assumption for now is that 1410 will keep up.

signal ADDR:      STD_LOGIC_VECTOR(13 downto 0);
signal LOAD_DATA: STD_LOGIC_VECTOR(7 downto 0);
signal DATA_LAST: STD_LOGIC := '0';

signal ADDR_COUNTER: INTEGER RANGE 0 to 3;

begin

loader_process: process(FPGA_CLK, RESET, loaderState, loaderAction,
   FIFO_READ_DATA_VALID, FIFO_EMPTY, FIFO_EMPTY_NEXT)

   begin

   if RESET = '1' then
      loaderState <= loader_RESET;
      loaderAction <= loader_Addr;

   elsif FPGA_CLK'event and FPGA_CLK = '1' then

      case loaderState is
      
         when loader_Reset => 
           DATA_LAST <= '0';
           ADDR_COUNTER <= 0;
           loaderState <= loader_WaitForChar;
           loaderAction <= loader_Addr;
            
         when loader_WaitForChar =>
            if(FIFO_EMPTY = '0') then
               FIFO_READ_ENABLE <= '1';
               loaderState <= loader_GetChar;
               loaderAction <= loaderAction;
            else
               loaderState <= loader_WaitForChar;
               loaderAction <= loaderAction;
            end if;
         
         when loader_GetChar =>
            if(FIFO_READ_DATA_VALID = '1') then

               case loaderAction is

                  when loader_Addr =>
                     if(FIFO_READ_DATA(6 downto 4) = MEMORY_LOADER_ADDRESS_MARK) then
                        -- Receiving address and see an address mark - OK
                        ADDR <= ADDR(8 downto 0) & FIFO_READ_DATA(3 downto 0);
                        if(ADDR_COUNTER = 3) then
                           loaderAction <= loader_Data;
                           DATA_LAST <= '0';
                           ADDR_COUNTER <= 0;
                        else
                           ADDR_COUNTER <= ADDR_COUNTER + 1;   
                           loaderAction <= loader_Addr;                     
                        end if;
                        loaderState <= loader_WaitForChar;
                     else 
                        -- Were not expecting an address mark...
                        loaderState <= loader_Reset;
                        loaderAction <= loader_Addr;
                     end if;

                  when loader_Data =>
                     if(FIFO_READ_DATA(6 downto 4) = MEMORY_LOADER_END_MARK) then
                        -- All Done
                        loaderState <= loader_Reset;
                        loaderAction <= loader_Addr; 
                     elsif((FIFO_READ_DATA(6 downto 4) = MEMORY_LOADER_DATA_0_MARK) AND 
                        (DATA_LAST = '0')) then
                        -- Received top bits of data...
                        LOAD_DATA(7 downto 4) <= FIFO_READ_DATA(3 downto 0);
                        DATA_LAST = '1';
                        loaderState <= loader_WaitForChar;
                        loaderAction <= loader_Data;
                     elsif((FIFO_READ_DATA(6 downto 4) = MEMORY_LOADER_DATA_1_MARK) AND
                        (DATA_LAST = '1')) then
                        -- Received bottom bits of data...
                        LOAD_DATA(3 downto 0) <= FIFO_READ_DATA(3 downto 0);
                        DATA_LAST = '0';
                        loaderState <= loader_Write;
                        loaderAction <= loader_Data;
                     else
                        --- ERROR
                        loaderState <= loader_Reset;
                        loaderAction <= loader_Addr;                        
                     end if;

                  end case;
                
               else
                  -- Should never actually get here...
                  loaderState <= loader_Reset;
                  loaderAction <= loader_addr;
               end if;  
             
            when loader_Write =>
               -- This can probably be combinatorial with "when" lists...
               loaderState <= loader_WrDone;
               loaderAction <= loader_Data;
               IBM1410_DIRECT_MEMORY_ADDRESS <= ADDR;
               IBM1410_DIRECT_MEMORY_WRITE_DATA <= LOAD_DATA;
               if(ADDR > '0111010100101111') then    -- 30000 and up
                  IBM1410_DIRECT_MEMORY_ENABLE = "1000";
                  IBM1410_DIRECT_MEMORY_WRITE_ENABLE = "1000";
               elsif(ADDR > '0100111000011111') then -- 20000 to 29999
                   IBM1410_DIRECT_MEMORY_ENABLE = "0100";
                   IBM1410_DIRECT_MEMORY_WRITE_ENABLE = "0100";
               elsif(ADDR > '0010011100001111') then -- 10000 to 19999
                   IBM1410_DIRECT_MEMORY_ENABLE = "0010";
                   IBM1410_DIRECT_MEMORY_WRITE_ENABLE = "0010";
               else                                  -- 00000 to 09999
                   IBM1410_DIRECT_MEMORY_ENABLE = "0001";
                   IBM1410_DIRECT_MEMORY_WRITE_ENABLE = "0001";
               endif;
               loaderState <= loader_WrDone;
               loaderAction <= loader_Addr;
                     
            when loader_WrDone =>
               IBM_DIRECT_MEMORY_ENABLE <= "0000";               
               IBM_DIRECT_MEMORY_WRITE_ENABLE <= "0000";
               loaderState <= loader_Getchar;
               loaderAction <= loader_Data;
            
      end case;
   
   end if;
   
   end process;

   -- Instantiate the FIFO ring buffer
   
   FIFO : ring_buffer
      generic map (
         RAM_WIDTH => MEMORY_LOADER_FIFO_WIDTH,
         RAM_DEPTH => MEMORY_LOADER_FIFO_SIZE
      )
      port map (
         clk => FPGA_CLK,
         rst => RESET,
         wr_en => SWITCH_FIFO_WRITE_ENABLE,
         wr_data => SWITCH_FIFO_WRITE_DATA,
         rd_en => FIFO_READ_ENABLE,
         rd_valid => FIFO_READ_DATA_VALID,
         rd_data => FIFO_READ_DATA,
         empty => FIFO_EMPTY,
         empty_next => FIFO_EMPTY_NEXT,
         full => FIFO_FULL,
         full_next => FIFO_FULL_NEXT,
         fill_count => OPEN
    );



end Behavioral;
